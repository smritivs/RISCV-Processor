module alu #(
    parameter DATA_WIDTH = 32)
