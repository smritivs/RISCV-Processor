module alu #(
    parameter DATA_WIDTH = 32
    )(
    input [DATA_WIDTH-1:0] a,b,
    input [5:0] alu_controls,
    input funct3b0,
    output reg [DATA_WIDTH-1:0] res
);

always @(*) begin
    case(alu_controls)
        6'b000000: res = a+b;
        6'b000001: res = a-b;
        6'b000010: res = a << (b[4:0]);
        6'b000011: res = ($signed(a) < $signed(b)) ? 32'd1 : 32'd0;
        6'b000100: res = ($unsigned(a) < $unsigned(b)) ? 32'd1 : 32'd0;
        6'b000101: res = a^b;
        6'b000110: res = a >> (b[4:0]);
        6'b000111: res = $signed(a) >>> (b[4:0]);
        6'b001000: res = a | b;
        6'b001001: res = a & b;
        6'b001010: res = ((a == b) ^ funct3b0) ? 32'd1 : 32'd0;
        6'b001011: res = ((a < b) ^ funct3b0) ? 32'd1 : 32'd0;
        6'b001100: res = (($signed(a) < $signed(b)) ^ funct3b0) ? 32'd1 : 32'd0;
        6'b001101: res = b;
        // p type
        6'b010000: res = {(a[31:16]+b[31:16]) << 16,a[15:0]+b[15:0]};
        6'b010001: res = {(a[31:16]-b[31:16]) << 16,a[15:0]-b[15:0]};
        6'b010010: res = {(a[31:16]+b[31:16]) << 16,a[15:0]-b[15:0]};
        6'b010011: res = {(a[31:16]-b[31:16]) << 16,a[15:0]+b[15:0]};
        6'b010100: res = {(a[31:24]+b[31:24]) << 24,(a[23:16]+b[23:16]) << 16,(a[15:8]+b[15:8]) << 8,a[7:0]+b[7:0]};
        6'b010101: res = {(a[31:24]-b[31:24]) << 24,(a[23:16]-b[23:16]) << 16,(a[15:8]-b[15:8]) << 8,a[7:0]-b[7:0]};
        6'b010110: res = {($signed(a[31:16]) >>> b[20:16]) << 16, $signed(a[15:0]) >> b[4:0]};
        6'b011000: res = {(a[31:16] >> b[20:16]) << 16, a[15:0] >> b[4:0]};
        6'b011010: res = {(a[31:16] << b[20:16]) << 16,a[15:0] << b[4:0]};
        6'b011100: res = {($signed(a[31:24]) >>> b[28:24]) << 24, ($signed(a[23:16]) >>> b[20:16]) << 16, ($signed(a[15:8]) >>> b[12:8]) << 8, $signed(a[7:0]) >>> b[4:0]};
        6'b011110: res = {((a[31:24]) >> b[28:24]) << 24, ((a[23:16]) >> b[20:16]) << 16, ((a[15:8]) >> b[12:8]) << 8, (a[7:0]) >> b[4:0]};
        6'b100000: res = {((a[31:24]) << b[28:24]) << 24, ((a[23:16]) << b[20:16]) << 16, ((a[15:8]) << b[12:8]) << 8, (a[7:0]) << b[4:0]};
        6'b100010: res = {($signed(a[31:16])*$signed(b[31:16])) << 16,$signed(a[15:0])+$signed(b[15:0])};
        6'b100011: res = {(a[31:16]*b[31:16]) << 16,a[15:0]*b[15:0]};
        6'b100100: res = {($signed(a[31:24])*$signed(b[31:24])) << 24,($signed(a[23:16])*$signed(b[23:16])) << 16,($signed(a[15:8])*$signed(b[15:8])) << 8,$signed(a[7:0])*$signed(b[7:0])};
        6'b100101: res = {(a[31:24]*b[31:24]) << 24,(a[23:16]*b[23:16]) << 16,(a[15:8]*b[15:8]) << 8,a[7:0]*b[7:0]};
        default: res = 32'd0;
    endcase
end
endmodule
