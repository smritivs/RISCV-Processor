module alu_decoder(
    input [2:0] alu_op
    );

endmodule
