module top()
// Instantiate various modules for linting purposes


endmodule